// Code your testbench here
// or browse Examples
`include "test_bench_new.sv"
//`include "test_bench2_new.sv"
//`include "test_bench3_new.sv"
// `include "Top.sv"
//`include "test0.txt"
//`include "test1.txt"
//`include "test2.txt"
//`include "test3.txt"
//`include "test4.txt"
//`include "test5.txt"
//`include "test6.txt"
//`include "test7.txt"
//`include "test8.txt"
//`include "test9.txt"
//`include "program1assembly.txt"