// Code your design here
`include "Top.sv"
`include "JLUT.sv"
`include "ProgCtr.sv"
`include "InstROM.sv"
`include "Ctrl.sv"
`include "RegFile.sv"
`include "ALU.sv"
`include "DMem.sv"
`include "ImmToRegMux.sv"
`include "MemToRegMux.sv"